module IDCT_tran();
endmodule
