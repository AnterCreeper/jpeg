module IDCT_mul();
endmodule
